module adder(
	
);



endmodule