module add_32(
	input [31:0] x, y,
	input C0,
	output C32,
	output [31:0] S
);
	
	wire G_0, P_0, G_1, P_1, G_2, P_2, G_3, P_3, G_4, P_4, G_5, P_5, G_6, P_6, G_7, P_7, C4, C8, C12, C16, C20, C24, C28;

	
	add_4 add_0_3(x[3:0], y[3:0], C0, S[3:0], G_0, P_0);
	
	add_4 add_4_7(x[7:4], y[7:4], C4, S[7:4], G_1, P_1);
	
	add_4 add_8_11(x[11:8], y[11:8], C8, S[11:8], G_2, P_2);
	
	add_4 add_12_15(x[15:12], y[15:12], C12, S[15:12], G_3, P_3);
	
	add_4 add_16_19(x[19:16], y[19:16], C16, S[19:16], G_4, P_4);
	
	add_4 add_20_23(x[23:20], y[23:20], C20, S[23:20], G_5, P_5);
	
	add_4 add_24_27(x[27:24], y[27:24], C24, S[27:24], G_6, P_6);
	
	add_4 add_28_31(x[31:28], y[31:28], C28, S[31:28], G_7, P_7);

	
	look_ahead_32 lk_32(
			C0, G_0, P_0, G_1, P_1, G_2, P_2, G_3, P_3, G_4, P_4, G_5, P_5, G_6, P_6, G_7, P_7, 
			C4, C8, C12, C16, C20, C24, C28, C32
	);
	

endmodule
