module look_ahead_16 (
	
);



endmodule
